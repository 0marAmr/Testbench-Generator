module FA_tb;

reg A, B, C_in;
wire S, C_out;

initial begin

end

endmodule